`include "base_seq_item.sv"
`include "rst_seq.sv"
`include "wr_seq.sv"
`include "base_seq.sv"
`include "base_seqr.sv"
`include "base_drv.sv"
`include "base_mon.sv"
`include "base_agt.sv"
`include "base_scb.sv"
`include "base_env.sv"
`include "base_test.sv"
