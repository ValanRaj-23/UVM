	`include "base_seq_item.sv"
	`include "rst_seq.sv"
	`include "write_seq.sv"
	`include "read_seq.sv"
	`include "base_seq.sv"
	`include "base_seqr.sv"
	`include "base_driver.sv"
	`include "base_monitor.sv"
	`include "base_scb.sv"
	`include "base_agent.sv"
	`include "base_env.sv"
	`include "base_test.sv"
